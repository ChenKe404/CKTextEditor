                
battle.ini       *   Brotherhood of Nod Campaign - Deus ex Kane    $   GDI Campaign - Evolutionary Response    mission.ini    J      A New Beginning    �  Another possible location of the Prototype Manufacturing Facility. Use the mutants to locate the position of the production facility. They must remain undetected. If Nod suspects enemy forces, they will cloak their production facility and deploy troops to destroy them. If the mutants can hide from the Nod troops for a short period, then Nod will assume the area is clear and uncloak the base. Once we record the location of the base, GDI Dropships will arrive with reinforcements.@@Objective One: Using Mutants you must locate the Prototype Manufacturing Facility.@@Objective Two: Once the facility is located reinforcements will be sent into help construct a base. You are to destroy the manufacturing facility at this time.    o  BE ADVISED: Kane is determined to destroy you. He knows the Kodiak cannot lift off during an ion storm and has chosen this moment to attack. The Kodiak must be protected until the storm abates. The storm will interfere with certain types of equipment so expect some malfunction.@@Objective One: Protect the Kodiak at all costs.@@Objective Two: Destroy all Nod forces.       Blackout       Capture Hammerfest Base       Capture Jake McNeil       Capture Train Station       Capture Umagon    �  Control of the mutants is in our grasp. Their headquarters is located to the north of your drop-off position. The units you will need to implicate GDI in this deception can be obtained by capturing the rest of the GDI base that you will start in. Do not mar the Brotherhoods name any further. Allow the blame to fall squarely upon Solomon's shoulders.@@Objective One: Capture the enemy Construction Yard awaiting you.@@Objective Two: Use GDI units to destroy the mutant's base.       Defend Crash Site       Destroy Chemical Missile Plant       Destroy Chemical Supply       Destroy GDI Research Facility       Destroy Mammoth Mk.II Prototype       Destroy Prototype Facility       Destroy Radar Array       Destroy Vega's Base       Destroy Vega's Dam    �   Destroy the three relay stations and the radar array to blackout Nod's sensor net. This will make rescuing Tratos easier, as Nod will not be as quick to detect you.@@Objective One: Destroy the three relay stations.@@Objective Two: Destroy the radar array.       Detroy Hassan's Temple    �  Emergency transmissions from GDI forces in this region indicate that Phoenix Base is under attack from Nod troops. It is imperative that the base be restored by building a Tiberium Refinery and a Barracks. Once the base is functional, all Nod forces in the area must be destroyed.@@Objective One: Build a Tiberium Refinery.@@Objective Two: Build a Barracks.@@Objective Three: Destroy all Nod forces.       Escort Bio-toxin Trucks       Establish Nod Presence       Eviction Notice       Final Conflict       Free Rebel Commander    �  GDI forces in this sector have found something unusual and large that crashed nearby. Nod has taken an intense interest in whatever it is, so naturally we are interested as well. Locate the object from the reports and capture any Nod Technology Centers in the area that might have uncovered clues as to the identity of the object.@@Objective One: Locate the Crash Site.@@Objective Two: Capture any Nod Technology Centers.    [  GDI has secured the Holy Ground the temple rests on. Your objective is simple, locate it and remove the GDI incursion. They are not expecting any Nod forces, so the element of surprise is yours. The temple and its knowledge must remain intact. One vision, One purpose!@@Object One: Locate the Temple of Nod.@@Objective Two: Destroy all GDI forces.    �  GDI has stored the firing codes for its Ion Cannon in three separate Comm centers. The centers are isolated in a valley and poorly guarded. We do not have the forces available for a full-scale assault. However, a small infiltration team led by the Chameleon Spy has a reasonable chance of success. Once the Spy has the codes, he must be evacuated safely.@@Objective One: Infiltrate the Comm centers and steal the codes.@@Objective Two: Evacuate the Chameleon Spy.      GDI is set to test the prototype of their new weapon, the Mammoth Mark II. It is vital that we sabotage their production of this monster as soon as possible. Before we can do that however, we need to know where the test is being held. Send a Chameleon Spy into one of the Radar Facilities. The coordinates to the testing ground should be stored there. Be careful of the patrols in the area - we have only one spy available. Once we have the location of the test, construct a base and destroy the prototype. You now have access to the new Banshee aircraft, which should prove useful. Destroying the remainder of the GDI base is at your discretion, but the Mammoth MUST be destroyed.@@Objective One: Spy on one of the GDI Comm Centers.@@Objective Two: Destroy the Mammoth Mark II prototype.    �  Hammerfest base has been overrun by Nod troops. The Firestorm walls block direct approach, so another route must be found back into the complex. Using hover MLRS and waterways for access, find a way back to the GDI base and re-capture it. Once the base is back in GDI hands, destroy all Nod forces in the area.@@Objective One: Find a way back to the GDI base.@@Objective Two: Re-capture the base with engineers.@@Objective Three: Destroy all Nod forces in the area.    =  Hassan is determined to stop you at any cost. He has pursued us back to a small base near his HQ. We must fend off his assault and build a Tiberium Refinery so we have the means to strike back.@@Objective One: Get production online by building a Tiberium Refinery.@@Objective Two: Destroy all of Hassan's Elite Guard.    �  Hassan spreads his propaganda to the Brotherhood through a nearby TV station. With the Brotherhood in chaos, the opportunity to divide Hassan from his followers presents itself. Capture the TV station and those once loyal to Kane's technology of peace will return to the fold. And as for Hassan's pathetic guards - crush them.@@Objective One: Capture the TV station to the east.@@Objective Two: Destroy Hassan's Elite Guard.    �  If the upcoming GDI attack on the missile sites is to succeed, C4 must be planted at all six power stations. The power grid is well protected, but the train should carry the demolition team and the mutants through the gates and past the guards. If Nod forces discover the demolition team and sound the alert, take out the power plants by any means available.@@Objective One: Plant C4 at the power plants.       Illegal Data Transfer    �  Impulses scanned from signatures emanating from Cairo suggest Kane will launch his world-altering missile within hours. You must destroy the Pyramid Temple before he has a chance to launch. There are no other strategies.@@Objective One: Clear the zone for MCV Dropship deployment.@@Objective Two: Destroy the ICBM launchers.@@Objective Three: Destroy the Pyramid Temple.@@Objective Four: Destroy all Nod forces.    �  In order for our ICBMs to shoot down the Philadelphia, they must be able to triangulate the station's position. Our spies have placed beacons at the optimal deployment locations. Once the launchers have been moved to the beacons, the station's fate is sealed and the Temple of Nod may be built. Move with all due haste. If the Philadelphia is able to complete three orbits, it will lock onto our position and destroy Kane's plans.@@Objective One: Deploy ICBM launchers at the three beacons.    ?  It is imperative that you prevent the train carrying the crystals from reaching the Nod base. Recent ice melts in the region have washed out the only train bridge. However, Nod engineers are on their way to repair it, so you must move quickly. If you can get to the train before the bridge is repaired, we can recover the crystals with little trouble. Otherwise, we will have to assault the Nod base to reclaim the crystals. Remember, to stop the train, you must destroy the locomotive, not the cars, but the cargo car holds the crystals.@@Objective One: Locate the train and destroy the locomotive before Nod engineers repair the bridge. The cargo car holds the crystals.@@Objective Two: If the bridge is repaired and the train successfully reaches the Nod base, then you must locate and destroy this base to recover the crystals.    -  Jake McNeil, brother of one of GDI's commanders, will be leading an inspection tour to a small GDI outpost in this area. His knowledge of GDI activities could be of great benefit to Nod's cause. Capture the GDI outpost with engineers, then disguise the base as GDI's and wait for Jake to make his inspection. When the signal is given, use the Toxin soldiers provided to "persuade" Jake to join Nod's forces. Once he is under our influence, EVAC him at the designated site.@@@Be very careful not to alert GDI until we are ready to strike. If they detect Nod forces in the area, they will surely try to evacuate Jake. If GDI is alerted, be sure to get to Jake before he can leave the area.@@Objective One: Capture the GDI outpost.@@Objective Two: Capture Jake.@@Objective Three: EVAC Jake at the specified location.       Mine Power Grid    �  Nod forces were recently forced out of this area. However, spies report that the Nod bio-toxin facility has not yet been destroyed by GDI troops. The Cyborg Commando and his team should be able to slip through the main GDI force and recover two tankers full of bio-toxin - provided we act quickly.@@Objective One: Locate the bio-toxin trucks.@@Objective Two: Escort the trucks to the checkpoint east of the base.    %  Nod has positioned a supply base in the area near a civilian train station. We can use the train and supplies to infiltrate the larger Nod base to the east. Avoiding patrols where possible and destroy all the Nod structures in the area. Once the area is secure, capture the train station for our use. DO NOT destroy the station or the train, as they are vital to our plans. Engineers and other reinforcements are available, but not unlimited - do not waste them.@@Objective One: Destroy all Nod structures.@@Objective Two: Capture the train station.    �  Nod is experimenting on mutant survivors at a facility in this sector. Among them is Tratos, leader of the mutants. Using Umagon's strike team, rescue Tratos from imprisonment and EVAC him at the specified site. Once complete, move in with GDI forces and destroy the Nod base and the prison test facility.@@Objective One: Rescue Tratos from prison.@@Objective Two: EVAC Tratos at specified site.@@Objective Three: Destroy the Nod base and test facility.    |  Nod's main chemical missile plant is located in this area. It is responsible for the large amount of Tiberium poisoning and accelerated mutations of wildlife in the surrounding areas. Destroying this facility will prevent Nod from furthering the acceleration of Tiberium poisoning on the planet.@@Objective One: Destroy Nod's missile silos.@@Objective Two: Destroy all Nod forces.    �  One of two possible locations of the Prototype Manufacturing Facility. Use the mutants to locate the position of the production facility. The mutants must remain undetected. If Nod suspects enemy forces in the area, they will cloak the facility and deploy troops to destroy them. If the mutants can hide from the Nod troops for a short period, the base will assume the area is clear and uncloak. Once we record the location of the base, GDI Dropships will arrive with reinforcements.@@Objective One: Using mutants you must locate the Prototype Manufacturing Facility.@@Objective Two: Once the facility is located, reinforcements will be sent in to help construct a base. You are to destroy the Manufacturing Facility at this time.       Protect Waste Convoys       Reinforce Phoenix Base       Rescue Prisoners       Rescue Tratos       Retaliation       Retrieve Disrupter Crystals       Salvage Operation       Secure Crash Site       Secure The Region       Sheep's Clothing    K  Taking out this weak position of GDI forces will allow us to reclaim our Sarajevo temple without interruption. Move in under the cover of an ion storm - while GDI's communications will be down. Take out the Radar Facility before the storm abates.@@Objective One: Locate and destroy the GDI Radar Facility before the ion storm ends.    �  The Cyborg Commando has been sent in to retrieve you. Once free, rendezvous with your rescue team to the south. Use them to locate and free Oxanna. She will soon be transported to the main GDI facility, optimal chances for success rely on obtaining her before she is transported. After she has been freed, commandeer a GDI transport to make your escape.@@Objective One: Locate and free Oxanna.@@Objective Two: Steal a GDI transport to make an escape.    K  The Infidel, Hassan, has been tracked to this region of Cairo. Build a base and eliminate this would-be pharaoh, the pretender to Kane's throne.@@Objective One: Cross the bridge and destroy the enemies on the far side.@@Objective Two: Deploy your MCV and begin building a base.@@Objective Three: Locate and destroy Hassan's Temple.       The Messiah Returns    �  The Nod base in this sector has been overrun by Tiberium life forms. Weedeaters have proven to be effective against the Tiberium creatures, but we must move reinforcements in quickly before the base is completely destroyed. Once the situation has been stabilized, the GDI base in the area must be eliminated.@@Objective One: Locate and secure the old base.@@Objective Two: Destroy the GDI base.    g  The Nod forces that attacked Phoenix Base have been traced back to a small base in this sector. Orders received from GDI Command state that the Nod base must be destroyed. However, there is a significant civilian population in the immediate area that must be evacuated by ORCA Transport before the fighting gets too heavy. Before the Transports can safely land, all seven SAM sites must be destroyed. Once the civilians have been evacuated, the Nod base can be destroyed.@@Objective One: Deploy the M.C.V. and begin building a base.@@Objective Two: Destroy all Nod SAM sites.@@Objective Three: Destroy the Nod base.    �  The alien craft is located in this region. FIND IT! The area is infested with GDI, so stealth would be to your advantage. Once the craft is located get an engineer inside to retrieve the Tacitus. And, should you encounter Vega's forces - consider them expendable.@@Objective One: Locate the crashed UFO and retrieve Kane's artifacts.@@Objective Two: Stop the transport of the Tacitus at all costs.    '  The hydroelectric dams in this area provide Vega's island fortress with almost limitless power. Destroying the dams will seriously cripple Vega's perimeter defenses and allow GDI to bring more weapons to bear against Vega's base.@@The dams are heavily fortified, so attacking them directly is not the best option. Surveillance indicates the key to destroying the dams lies in the destruction of two regulator stations. Without them, the dams' generators will overload and the dams will self destruct.@@Objective One: Destroy the dams any way possible.    U  The mutant female may be trying to reach the underground railway system located in New Detroit. Move in and control the station before she arrives. If she boards the train then it must be stopped. This may be our last chance at capturing the abomination.@@Objective One: Locate the train station in the area and capture it before Umagon flies in and boards the train to escape into the underground.@Objective Two: If Umagon boards the train before you have captured the station then you must stop the train before it leaves the region. Destroy the locomotive and we will be able to capture Umagon.    �  The research facility in this sector must be destroyed before the GDI scientists perfect their Tiberium reduction technology. If Nod forces are to establish a base in the area, the GDI patrols must be eliminated. The mutants may prove to be useful allies.@@Objective One: Contact the mutants@@Objective Two: Clear GDI forces away from the tunnel and main road.@@Objective Three: Locate the research facility.@Objective Four: Destroy the research facility.    �  The road through this sector is a vital supply link. If a foothold is firmly established and a Tiberium Waste Facility is built, Nod chemical missiles can be launched from the region. The GDI base in the area has no defense against the missiles, and can be destroyed at your leisure once the waste convoys start arriving.@@Objective One: Establish a base and build a Tiberium Waste Facility@@Objective Two: Destroy the GDI base.    /  This chemical supply station is providing vast quantities of Tiberium toxins to a number of Nod research programs in the area. Destroying this site will seriously hinder further Nod research, and prevent this base from transporting reinforcements to others in the sector.@@Intelligence reports advise caution when near any of the chemical tanks and facilities, as the toxins contained within are highly corrosive and equally deadly to soldiers and vehicles.@@Objective One: Find a suitable location for a base. Objective Two: Destroy the Nod Chemical station.    �  Umagon has requested help to rescue her people from a Nod prison. The prison is located on an island to the east. Nod has a strong force in the area, both in outposts and spread through the nearby city. We have limited resources and no reinforcements are available, so avoiding patrols is vital to your success. Umagon has a team in the area already - if you can find them, they may assist you. Make your way to the prison and release the hostages. Once the prison is secure, we will send a transport to evacuate Umagon's people. There may be SAM sites nearby, so make sure the way is clear for the transport.@@Objective One: Locate the Nod prison.@@Objective Two: Release and evacuate the prisoners.    �  Vega's base of operations is in the area. It is heavily guarded by SAM sites, and a secondary outpost provides reinforcements. Destroy all Nod forces in the area, but capture Vega's Pyramid intact - there is information there that we can use. You will have only limited troops until the SAM sites are neutralized one way or another.@@Objective One: Destroy the Nod base.@@Objective Two: Capture Vega's Pyramid.       Villainess in Distress    8  We have become aware of an imprisoned commander in this region who WAS loyal to Hassan. Free him and his forces and they should be sympathetic to our cause - and help in the capture of Hassan. The commander may have information vital to Hassan's movement.@@Objective One: Locate and free the Rebel Nod Commander.       Weather the Storm      Whatever is contained in this craft, it is apparent that Nod doesn't want GDI to have it. Protect the crashed UFO until GDI reinforcements can arrive to fortify the area.@@Objective One: Survive until reinforcements can arrive.@@Objective Two: Prevent Nod from destroying the UFO.    E  You must reach the medical colony in the region without being prematurely detected by GDI and forcing a base evacuation. To prevent this, consider first destroying the three sensor towers protecting the base. Our new artillery unit should be sufficient for the job. Once inside the base, the capture of the mutant female should be easy.@@Objective One: Find and destroy the GDI sensor towers without getting too close and getting detected by them.@@Objective Two: Once the towers are destroyed, move on the base and capture the medical colony before Umagon, the Mutant, can escape.    	rules.ini         2nd National Bank       Abandoned Factory       Abandoned Warehouse       Abandoned Wharehouse       Adam's House       Adult Visceroid       Advanced Power Plant       Alex-gators petshop just ahead!       Alkaline's Battery Superstore       AlphaLightPost       Ambrose Lounge       Ammo Crates       Amphibious APC       Archer Asylum    	   Artillery       Attack Buggy       Attack Cycle    
   Automobile       Baby Visceroid       Banshee       Barracks       Billy Bob's Harvester school       Blue Light Post       Bostic Tower       Boxes       Bridge 1       Bridge 2       Bridge repair hut       Business Offices    	   Cargo Car       Carryall       Chameleon Spy       Chem Spray Infantry       Chemical Missile       Church    	   City Hall       Civilian       Civilian Armory       Civilian Array       Civilian Hospital       Clear Rock #1       Clear Rock #2       Clear Rock #3       Clear Rock #4       Clear Rock #5       Component Tower       Concrete Wall       Connelly Court Apts.       Construction Yard       Crash 1       Crash 2       Crash 3       Crash 4       Crash 5       Crate       Cyborg       Cyborg Commando       Daily Sun Times       Dam       Deluxe Accomodations       Denzil's Last Chance Motel       Deployed Artillery       Deployed ICBM       Deployed Sensor Array       Deployed Tick Tank       Devil's Tongue       Disc Thrower    	   Disruptor       Disruptor Turret       Drink YEO-CA Cola!       Drop Pod       Dropship       Drum    
   E.M. Pulse    
   EMP Cannon       Eat at Rade's Roadhouse       Energy Transformer       Engineer       Ferbie's 4 Sale       Field Generator       Fill'er Up-Pump'N'Go       Fire Storm Generator       Firestorm Defense       Firestorm Wall Section       Flying Gas Tank       Flying Tire       GDI       GDI Hunter-Seeker    
   GDI Kodiak       GDI Power Plant       GDI Tech Center       GDI Upgrade Center       GDI War Factory       Gas Pump    	   Gas Pumps       Gas Station       Gas Station Sign       Gate       Ghost Stalker       Goodie Crate       Green Building       Green Light Post    
   Greenhouse       Hamburgers $.99       Hand Of Nod       Harpy    	   Harvester       Helipad       Hewitt Hair Salon       Highrise Hotel    
   Hover MLRS       Hunter Seeker       Hunting Lodge       Ice Floe       Invisible Blue Light Post       Invisible Green Light Post       Invisible Light Post       Invisible Purple Light Post       Invisible Red Light Post       Invisible Yellow Light Post    
   Ion Cannon       Ion Cannon Uplink       JP       Join GDI: We save lives.       Jumpjet Infantry       Kaspm's Tiberium Warhouse       Kettler's Place       Large Tiberium       Laser       Laser Fence Post       Laser Fence Section       Leary Traveller Inn       Light Infantry    
   Light Post       Light Tower       Lightner's Luxury Suites       Local Inn & Lodging       Local Store    
   Locomotive       Long's Home    
   Low Bridge       Low Bridge End 1       Low Bridge End 2       Low Bridge End 3       Low Bridge End 4       Mammoth Mk.II       Mammoth Tank       Mammoth Tank Turret       Medic       Meteorite01       Meteorite02       Miele Manor       Missile Launcher       Missile Silo       Mobile Construction Vehicle       Mobile Repair Vehicle       Mobile Sensor Array       Multi-Missile       Mutant       Mutant Hijacker       Mutant Sergeant       Mutant Soldier       NOD       NOD Montauk       NOD Power Plant       NOD Pyramid    	   NOD Radar       NOD Tech Center       Negative Light Post       Negative Red Light       No escape from Archer's Asylum!       Nod Hunter-Seeker       Nod Wall       Nod War Factory       Obelisk of Light       Observation Tower       Office Building       Old Advanced Power Plant       Old Construction Yard       Old Refinery    	   Old Silos    
   Old Temple       Old Weapons Factory       Only 11 miles to Zydeko's cafe!       Orange Light Post       Orca Bomber       Orca Fighter       Orca Transport       Oxanna       Palette       Pannullo's hacienda es bueno       Panullo Hacienda       Pavement       Pickup Truck       Port-A-Shack       Port-A-Shack Deluxe       Power Turbine       Purple Light Post       Pyramid       RPG Upgrade       Radar       Rade's Roadhouse       Railroad Bridge 1       Railroad Bridge 2       Recreational Vehicle       Red Light Post       Rocket Infantry       Rooms $29 a nite       SAM Upgrade       Sam       Sand Rock #1       Sand Rock #2       Sand Rock #3       Sand Rock #4       Sand Rock #5       Sandbags       Sandberg and Son's    
   School Bus       Scrap Metal Debris    
   Scrin Ship       Seeker Control       Service Depot       Slavick       Solar Panel       Stealth Generator       Stealth Tank       Stop in at Hewitt's hair salon       Subterranean APC       Subterranean Dwelling       TacticX games rock!       Tall's Residence    
   Technician       Temp Housing       Temple of NOD       The Projects       Threat Rating Node       Tiberian Fiend    ,   Tiberian Sun -- Official Rules of Engagement       Tiberium       Tiberium (Blue)       Tiberium (Green)       Tiberium (Large)       Tiberium Aboreus       Tiberium Cruentus       Tiberium Refinery       Tiberium Riparius       Tiberium Silo       Tiberium Tree       Tiberium Veins       Tiberium Vinifera       Tiberium Waste Facility       TiberiumCrystal01       TiberiumCrystal02       TiberiumShard    	   Tick Tank       Titan       Track EW       Track NS    
   Track NeSw    
   Track NwSe    	   Train Car       Train Tracks       Tratos       Tree       Truck       Truck (loaded)       Umagon       Urban Housing       Urban Storefront       Vega's Pyramid       Veinhole Monster       Veinhole Monster Dummy       Veinhole Tree       Visit Scenic Las Vegas       Vulcan Cannon       WS Logging Company       WW Surf and Turf hits the spot!       Water Purifier    
   Water Tank    
   Waystation    
   Weed Eater       Westwood Stock Exchange    	   Wolverine       YEO-CA Cola Corp.       Yee's Discount Liquor       Yellow Light Post    tutorial.ini    �      ****BROADCASTING****       1...       2,       Alert! GDI presence detected!        Alert! Prison break in progress!       BATTLEFIELD CONTROL ESTABLISHED    !   Base perimeter has been breached!    2   Beware Tiberium is lethal to unprotected infantry.    '   Build more infantry to defend the base!       Bullet train departing.    �   CABAL: During the Ion Storm their Radar/Communications will be down. Now is the opportune time to hit them before the storm abates.    ]   CABAL: Establish a foothold on the far side of this bridge and an MCV will be sent in to you.    �   CABAL: Find and capture the train station before Umagon arrives. If she manages to make it onto a train then destroy it before she can escape.    2   CABAL: GDI Communications have been reestablished.    B   CABAL: General Vega, the generators are online.  SAM sites active.    M   CABAL: General Vega, the secondary generators will come online in 20 minutes.    :   CABAL: Hassan's Base has been alerted. Attack is imminent.    (   CABAL: MCV has arrived to the southeast.    .   CABAL: Philadelphia orbit tracking commencing!    #   CABAL: Slavik lost, mission failed.    S   CABAL: With the train destroyed Umagon will be stranded.  Find her and capture her.       CAUTION: THIN ICE.    W   Captured Commander: All right! Now get me to your drop-off site and into the evac unit.       Civilian city is under attack!    .   Clear the zone for M.C.V. dropship deployment!       Codes located.       Convoy destroyed.    ;   Current weapon range insufficient. Weapon drop in progress.    7   Deploy the M.C.V. by double left clicking on the M.C.V.    H   Destroy the 7 SAM sites on the ridge to clear the way for our dropships.       Detonate C4 when ready.       Down with Hassan!!!    +   ESTABLISHING BATTLEFIELD CONTROL - Standby!    j   EVA: Alert! The bridge has been fixed and the Nod train is moving to its final destination within the base    [   EVA: GDI reinforcements have arrived. Mammoth Mk II enroute.  Estimated ETA in 2 minutes...    %   EVA: Ghostalker lost, mission failed.       EVA: Mammoth Mk II has arrived.    !   EVA: Mcneil lost, mission failed.    ^   EVA: Penetrate their base, destroy that cargo car and retrieve the crate holding the crystals.    `   EVA: The bridge has been repaired and the train is making it's way to the Nod base in the south.    X   EVA: The cargo car of that train contains the crate of crystals that you are to recover.    8   EVA: The crystals have been retrieved, mission complete.    !   EVA: Umagon lost, mission failed.    l   EVA: We are currently tracking the Nod train carrying the target cargo.  Intel states that the bridge is out    "   Eye of the storm has been entered.        Firestorm perimeter deactivated.       First launcher deployed.    /   GDI Forces Spotted! Falling back to alert base.    H   GDI Soldier: Shit, We're outnumbered! Return to base now and alert them.       GDI bullet train arriving.       GDI bullet train departing.       GDI dropship detected.    $   GDI forces spotted. Blow the bridge!       GDI has detected you.    ?   GDI is going after our extraction APC It must not be destroyed!    *   GDI: Hurry Jake! They're right behind you!    +   GDI: Jake, it's a trap! Get to the airbase!    6   GDI: Jake, it's good to see...Hey! What are you doing?    A   GDI: Jake, the transport will take 30 minutes to arrive. Hold on!    6   GDI: Now watch the effectiveness against ground units.    4   GDI: Patrol to base! Nod troops in area! Abort tour!    5   GDI: The MM2 is equally deadly to air-based assaults.    3   GDI: The MM2 is quite effective against structures.    6   GDI: This concludes the Mammoth Mark II demonstration.    G   GDI: We've lost the beacon. Extraction time will be delayed 15 minutes.    M   Ghost Stalker: If you can get me onto that train, we can do some real damage!    "   Harvest the Tiberium to the north.       Hassan Soldier: Hold them here!    )   Hey! Where'd all those shiners come from?    :   Hey... over here! Help... Destroy these trucks to free us.    +   Holy $#!+ its Nod! I have to warn the base.       ICBM destroyed!       ICBM launch detected.    +   ICBMs destroyed! Philidephia out of danger.    U   If your Tiberium Refinery is full, build Tiberium Silos to store the excess Tiberium.       Kodiak destroyed!       Kodiak in critical condition!       Kodiak under attack!       Laser Turrets! RUN FOR IT!       Launcher destroyed.    9   Looks like they're going to ship it out via bullet train.    5   Maximum efficiency for equipment can now be achieved.       Mission failed.    !   Move quickly, before they see us.       Mutant vermin detected.    P   Mutants: Damn, their base has been cloaked. We must wait for them to uncloak it.    5   Mutants: Hold a moment, while their fighters pass by.    @   Mutants: Liars! GDI is trying to help us! You will die for this!       Mutants: Okay, Go now.    N   Mutants: The charges are placed. We can get the laser wall down in 30 minutes.    d   Mutants: The production facility has been located. Send in the reinforcements and let's finish this.    4   Mutants: The wall is down - you are clear to attack!    D   New Objective: Get Ghost Stalker onto the train. Ghost must not die!    A   New secondary objective: Destroy primary AND secondary Nod bases.    8   Nod ICBMs detected. To stop them, DESTROY the launchers.    f   Nod base is heavily guarded by lasers. Suggestion: destroying power plants to west may cause overload.    X   Nod:  We can use these old units to our advantage.  Rerouting their control to you in 3,    I   Nod: All sensor arrays are down. Full area map generation dowloading now.    W   Nod: Commander, you have been provided with a direct satellite uplink for this mission.    ]   Nod: Look to your radar now and you will see the three locations of the mobile sensor arrays.    8   Nod: Umagon has been detected in the northeast quadrant.    1   Nod: Umagon has escaped. Your mission has failed.    Z   Nod: Umagon has reached the GDI base and is moving to board the train leaving this region.    b   Nod: Umagon is moving to board the northern train which leaves the region. Her escape is imminent.    [   Nod: Umagon's dropship transport has arrived and she is moving to board the southern train.    P   Nod: Umagon's dropship transport has been located and will arrive in 10 minutes.    9   Nod: Umagon's dropship transport will arrive in 1 minute.    :   Nod: Umagon's dropship transport will arrive in 5 minutes.    P   Note that your power is getting low. To get more power, build more Power Plants.    [   Now get an engineer over here to fix this bridge and I will alert Hassan to their presence.       O.K.! You're clear to enter.       Objective 1 complete.    Z   Objective 1: Build a Tiberium Refinery and begin harvesting the Tiberium to the southeast.    7   Objective 1: Capture Hassan's T.V. station to the east.    8   Objective 1: Capture the GDI base before McNeil arrives.    f   Objective 1: Capture the remaining GDI structures within this base to build a force to capture Tratos.    I   Objective 1: Contact the mutants - try searching near the local hospital.    8   Objective 1: Deploy the ICBM launchers near the beacons.    )   Objective 1: Destroy Nod missile complex.    (   Objective 1: Destroy all Nod structures.    7   Objective 1: Destroy all chemical missile launch sites.    1   Objective 1: Destroy all of Hassan's elite guard.    ,   Objective 1: Destroy all the chemical tanks.    %   Objective 1: Destroy the supply base.    B   Objective 1: Establish a base and build a Tiberium Waste Facility.       Objective 1: Establish a base.    $   Objective 1: Find and rescue Oxanna.    >   Objective 1: Infiltrate the GDI Communication Upgrade Centers.    )   Objective 1: Locate and free the mutants.    .   Objective 1: Locate and secure the crash site.    8   Objective 1: Locate the abandoned Nod base to the north.    N   Objective 1: Locate the crashed UFO and retrieve Kane's artifacts from inside.    *   Objective 1: Locate the old Temple of Nod.    %   Objective 1: Locate the toxin trucks.    2   Objective 1: Plant C4 on all ten Nod power plants.    -   Objective 1: Protect the Kodiak at all costs.    3   Objective 1: Remove all Nod presence from the area.    N   Objective 1: Spy on GDI comm center to learn the location of the weapons test.    5   Objective 1: Stop the launch of the Tiberium Missile.       Objective 2 complete.    6   Objective 2: Build a Barracks to create more infantry.    %   Objective 2: Build the Temple of Nod.    +   Objective 2: Capture Nod Technology Center.    $   Objective 2: Capture Vega's Pyramid.    :   Objective 2: Capture the train station. DO NOT DESTROY IT!    7   Objective 2: Clear both ends of the tunnel to the west.    .   Objective 2: Commandeer a transport to escape.    /   Objective 2: Destroy Hassan's elite guard base.    $   Objective 2: Destroy all Nod forces.    ,   Objective 2: Destroy all five Nod SAM sites.    "   Objective 2: Destroy the GDI base.    ;   Objective 2: Destroy the ICBMs targeted at the Philidephia.    3   Objective 2: Destroy the Mammoth Mark II prototype.    "   Objective 2: Destroy the Nod base.    I   Objective 2: Escort the toxin trucks past the GDI checkpoint to the east.    (   Objective 2: Evacuate the Chameleon Spy.    "   Objective 2: Evacuate the mutants.    �   Objective 2: Now find the Mutant Headquarters and knock on their door (attack it!). This should convince Tratos to be sympathetic to our cause.    (   Objective 2: Remove the GDI trespassers.    /   Objective 2: Retrieve the cargo from the train.    @   Objective 2: To get production online build a Tiberium Refinery.    @   Objective 2: Use Toxin Soldiers to "convince" McNeil to join us.    0   Objective 3: Destroy all Nod forces in the area.    $   Objective 3: Destroy all Nod forces.    =   Objective 3: Get McNeil into the APC at the extraction point.    7   Objective 3: Locate the research facility to the north.    +   Objective 4: Destroy the research facility.    '   Objective Reached: Civilians evacuated.    !   Objective Reached: Mutants freed.       Objective Reached: Site secure    .   Objective Reached: Technology Center captured.    7   Objective: Rescue captives from the prison to the east.       One launcher remaining.    F   Orca Transport: Negative on extraction until SAM sites are eliminated!    9   Our cover is blown! Capture McNeil by any means possible!    +   Oxanna is being moved to the main GDI base.       Oxanna located.       PEACE THROUGH POWER!    %   Perimeter secure. Deactivating alarm.       Philidelphia in range.    2   Power levels are low. Construct more Power Plants.       Power overload in progress...    :   Prevent the train from departing and retreive the Tacitus.    1   Proceed to the next Communication Upgrade Center.    *   Proceed with Tiberium Missile destruction.       Pull over for inspection!    )   Reentering ion storm, caution is advised.       SCROOGE!       STOP THAT TRAIN!       Second launcher deployed.    <   She is boarding a train bound for the GDI base in the south.    M   Sir! I believe there is an old GDI base near. It could be worth looking into.    8   Sir! The Tacitus is gone. Vega's men must've grabbed it.    p   Solomon: Change of plans - We have verified Vega's presence in the pyramid. CAPTURE the pyramid with Vega alive.    *   Sound the Alarm! Slavik's Forces are here!       Special objective complete.    0   Stand and Identify yourself in the name of Kane.        Stand forward and be recognized!    1   Stop! Don't Shoot! I was forced to work for them.    -   Storm abating. Commence attack on Nod forces.       Supplies found.       Tacitus has been acquired.    @   Take out this sentry post and I will show you their nearby base.       Thanks for the help!    ;   Thanks! We can use the supplies.  I'll go gather my people.    $   The Philadelphia has been destroyed!    %   The Philidelphia has left ICBM range.    .   The Philidelphia is passing within ICBM Range.       The Temple is under attack!    @   The temple has been discovered, NOW DESTROY the GDI trespassers.    ,   The traitors are coming, destroy the bridge!    0   They are sending a transmission to Sarajevo now.    ,   Third launcher deployed. Objective complete.       This map is under redesign.       Tiberium Missile launched.       Tiberium lifeform detected.    "   Tiberium waste convoy approaching.    A   To build or train left-click on the icons located in the sidebar.    V   To deploy a vehicle select it, place the cursor over the vehicle and left-click on it.    N   To repair a bridge, send an engineer into the repair hut near the bridge base.    c   To repair a structure left-click on the wrench icon in the sidebar and left-click on the structure.       Transport has arrived.       Transport lost.    ;   Tratos: Fight them my children, for the fate of our people.    V   Tratos: You have killed enough of my children, take me and be done with this violence.       Two launchers remaining.       UFO crash sight located.       Umagon: My people are nearby.    5   Umagon: My people are waiting somewhere to the north.    6   Use the Weedeater units to harvest the Tiberium veins.    1   Warning: Mission critical structure under attack.    ,   Warning: Mission critical unit under attack.    X   We have Hassan pinned and ready to be brought in Commander Slavick. Orders are complete.    *   We have to get this to Tratos immediately.    7   We should rendezvous with the rescue team to the south.       We will help.    ^   We've been touched by the spirit hand of Kane, and are ready to serve the technology of peace.    ?   What's the E.T.A. on that M.C.V.? This UFO gives me the creeps.    d   You have been provided with 2 Artillery units. Good hunting, reinforcements will be arriving soon...    =   Your venture has been quite unsuccessful, to state the least.    7   and we may hit the train before they repair the bridge.    C   to the South. Penetrate the bases defenses and retrieve that cargo.    